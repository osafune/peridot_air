// c4e_dvp_core_uart_to_avmm_bridge.v

// Generated using ACDS version 20.1 720

`timescale 1 ps / 1 ps
module c4e_dvp_core_uart_to_avmm_bridge (
		output wire [31:0] avm_address,       //   avm.address
		input  wire [31:0] avm_readdata,      //      .readdata
		output wire        avm_read,          //      .read
		output wire        avm_write,         //      .write
		output wire [31:0] avm_writedata,     //      .writedata
		input  wire        avm_waitrequest,   //      .waitrequest
		input  wire        avm_readdatavalid, //      .readdatavalid
		output wire [3:0]  avm_byteenable,    //      .byteenable
		input  wire        clk_clk,           //   clk.clk
		input  wire        reset_reset_n,     // reset.reset_n
		output wire        uart_txd,          //  uart.txd
		input  wire        uart_rxd,          //      .rxd
		input  wire        uart_cts,          //      .cts
		output wire        uart_rts           //      .rts
	);

	wire        sc_fifo_0_out_valid;                                    // sc_fifo_0:out_valid -> st_bytes_to_packets_0:in_valid
	wire  [7:0] sc_fifo_0_out_data;                                     // sc_fifo_0:out_data -> st_bytes_to_packets_0:in_data
	wire        sc_fifo_0_out_ready;                                    // st_bytes_to_packets_0:in_ready -> sc_fifo_0:out_ready
	wire        st_packets_to_bytes_0_out_bytes_stream_valid;           // st_packets_to_bytes_0:out_valid -> uart_to_bytes_0:in_valid
	wire  [7:0] st_packets_to_bytes_0_out_bytes_stream_data;            // st_packets_to_bytes_0:out_data -> uart_to_bytes_0:in_data
	wire        st_packets_to_bytes_0_out_bytes_stream_ready;           // uart_to_bytes_0:in_ready -> st_packets_to_bytes_0:out_ready
	wire        uart_to_bytes_0_source_valid;                           // uart_to_bytes_0:out_valid -> sc_fifo_0:in_valid
	wire  [7:0] uart_to_bytes_0_source_data;                            // uart_to_bytes_0:out_data -> sc_fifo_0:in_data
	wire        uart_to_bytes_0_source_ready;                           // sc_fifo_0:in_ready -> uart_to_bytes_0:out_ready
	wire        st_bytes_to_packets_0_out_packets_stream_valid;         // st_bytes_to_packets_0:out_valid -> avalon_st_adapter:in_0_valid
	wire  [7:0] st_bytes_to_packets_0_out_packets_stream_data;          // st_bytes_to_packets_0:out_data -> avalon_st_adapter:in_0_data
	wire        st_bytes_to_packets_0_out_packets_stream_ready;         // avalon_st_adapter:in_0_ready -> st_bytes_to_packets_0:out_ready
	wire  [7:0] st_bytes_to_packets_0_out_packets_stream_channel;       // st_bytes_to_packets_0:out_channel -> avalon_st_adapter:in_0_channel
	wire        st_bytes_to_packets_0_out_packets_stream_startofpacket; // st_bytes_to_packets_0:out_startofpacket -> avalon_st_adapter:in_0_startofpacket
	wire        st_bytes_to_packets_0_out_packets_stream_endofpacket;   // st_bytes_to_packets_0:out_endofpacket -> avalon_st_adapter:in_0_endofpacket
	wire        avalon_st_adapter_out_0_valid;                          // avalon_st_adapter:out_0_valid -> packets_to_master_0:in_valid
	wire  [7:0] avalon_st_adapter_out_0_data;                           // avalon_st_adapter:out_0_data -> packets_to_master_0:in_data
	wire        avalon_st_adapter_out_0_ready;                          // packets_to_master_0:in_ready -> avalon_st_adapter:out_0_ready
	wire        avalon_st_adapter_out_0_startofpacket;                  // avalon_st_adapter:out_0_startofpacket -> packets_to_master_0:in_startofpacket
	wire        avalon_st_adapter_out_0_endofpacket;                    // avalon_st_adapter:out_0_endofpacket -> packets_to_master_0:in_endofpacket
	wire        packets_to_master_0_out_stream_valid;                   // packets_to_master_0:out_valid -> avalon_st_adapter_001:in_0_valid
	wire  [7:0] packets_to_master_0_out_stream_data;                    // packets_to_master_0:out_data -> avalon_st_adapter_001:in_0_data
	wire        packets_to_master_0_out_stream_ready;                   // avalon_st_adapter_001:in_0_ready -> packets_to_master_0:out_ready
	wire        packets_to_master_0_out_stream_startofpacket;           // packets_to_master_0:out_startofpacket -> avalon_st_adapter_001:in_0_startofpacket
	wire        packets_to_master_0_out_stream_endofpacket;             // packets_to_master_0:out_endofpacket -> avalon_st_adapter_001:in_0_endofpacket
	wire        avalon_st_adapter_001_out_0_valid;                      // avalon_st_adapter_001:out_0_valid -> st_packets_to_bytes_0:in_valid
	wire  [7:0] avalon_st_adapter_001_out_0_data;                       // avalon_st_adapter_001:out_0_data -> st_packets_to_bytes_0:in_data
	wire        avalon_st_adapter_001_out_0_ready;                      // st_packets_to_bytes_0:in_ready -> avalon_st_adapter_001:out_0_ready
	wire  [7:0] avalon_st_adapter_001_out_0_channel;                    // avalon_st_adapter_001:out_0_channel -> st_packets_to_bytes_0:in_channel
	wire        avalon_st_adapter_001_out_0_startofpacket;              // avalon_st_adapter_001:out_0_startofpacket -> st_packets_to_bytes_0:in_startofpacket
	wire        avalon_st_adapter_001_out_0_endofpacket;                // avalon_st_adapter_001:out_0_endofpacket -> st_packets_to_bytes_0:in_endofpacket

	altera_avalon_packets_to_master #(
		.FAST_VER    (0),
		.FIFO_DEPTHS (2),
		.FIFO_WIDTHU (1)
	) packets_to_master_0 (
		.clk               (clk_clk),                                      //           clk.clk
		.reset_n           (reset_reset_n),                                //     clk_reset.reset_n
		.out_ready         (packets_to_master_0_out_stream_ready),         //    out_stream.ready
		.out_valid         (packets_to_master_0_out_stream_valid),         //              .valid
		.out_data          (packets_to_master_0_out_stream_data),          //              .data
		.out_startofpacket (packets_to_master_0_out_stream_startofpacket), //              .startofpacket
		.out_endofpacket   (packets_to_master_0_out_stream_endofpacket),   //              .endofpacket
		.in_ready          (avalon_st_adapter_out_0_ready),                //     in_stream.ready
		.in_valid          (avalon_st_adapter_out_0_valid),                //              .valid
		.in_data           (avalon_st_adapter_out_0_data),                 //              .data
		.in_startofpacket  (avalon_st_adapter_out_0_startofpacket),        //              .startofpacket
		.in_endofpacket    (avalon_st_adapter_out_0_endofpacket),          //              .endofpacket
		.address           (avm_address),                                  // avalon_master.address
		.readdata          (avm_readdata),                                 //              .readdata
		.read              (avm_read),                                     //              .read
		.write             (avm_write),                                    //              .write
		.writedata         (avm_writedata),                                //              .writedata
		.waitrequest       (avm_waitrequest),                              //              .waitrequest
		.readdatavalid     (avm_readdatavalid),                            //              .readdatavalid
		.byteenable        (avm_byteenable)                                //              .byteenable
	);

	altera_avalon_sc_fifo #(
		.SYMBOLS_PER_BEAT    (1),
		.BITS_PER_SYMBOL     (8),
		.FIFO_DEPTH          (256),
		.CHANNEL_WIDTH       (0),
		.ERROR_WIDTH         (0),
		.USE_PACKETS         (0),
		.USE_FILL_LEVEL      (0),
		.EMPTY_LATENCY       (3),
		.USE_MEMORY_BLOCKS   (1),
		.USE_STORE_FORWARD   (0),
		.USE_ALMOST_FULL_IF  (0),
		.USE_ALMOST_EMPTY_IF (0)
	) sc_fifo_0 (
		.clk               (clk_clk),                              //       clk.clk
		.reset             (~reset_reset_n),                       // clk_reset.reset
		.in_data           (uart_to_bytes_0_source_data),          //        in.data
		.in_valid          (uart_to_bytes_0_source_valid),         //          .valid
		.in_ready          (uart_to_bytes_0_source_ready),         //          .ready
		.out_data          (sc_fifo_0_out_data),                   //       out.data
		.out_valid         (sc_fifo_0_out_valid),                  //          .valid
		.out_ready         (sc_fifo_0_out_ready),                  //          .ready
		.csr_address       (2'b00),                                // (terminated)
		.csr_read          (1'b0),                                 // (terminated)
		.csr_write         (1'b0),                                 // (terminated)
		.csr_readdata      (),                                     // (terminated)
		.csr_writedata     (32'b00000000000000000000000000000000), // (terminated)
		.almost_full_data  (),                                     // (terminated)
		.almost_empty_data (),                                     // (terminated)
		.in_startofpacket  (1'b0),                                 // (terminated)
		.in_endofpacket    (1'b0),                                 // (terminated)
		.out_startofpacket (),                                     // (terminated)
		.out_endofpacket   (),                                     // (terminated)
		.in_empty          (1'b0),                                 // (terminated)
		.out_empty         (),                                     // (terminated)
		.in_error          (1'b0),                                 // (terminated)
		.out_error         (),                                     // (terminated)
		.in_channel        (1'b0),                                 // (terminated)
		.out_channel       ()                                      // (terminated)
	);

	altera_avalon_st_bytes_to_packets #(
		.CHANNEL_WIDTH (8),
		.ENCODING      (0)
	) st_bytes_to_packets_0 (
		.clk               (clk_clk),                                                //                clk.clk
		.reset_n           (reset_reset_n),                                          //          clk_reset.reset_n
		.out_channel       (st_bytes_to_packets_0_out_packets_stream_channel),       // out_packets_stream.channel
		.out_ready         (st_bytes_to_packets_0_out_packets_stream_ready),         //                   .ready
		.out_valid         (st_bytes_to_packets_0_out_packets_stream_valid),         //                   .valid
		.out_data          (st_bytes_to_packets_0_out_packets_stream_data),          //                   .data
		.out_startofpacket (st_bytes_to_packets_0_out_packets_stream_startofpacket), //                   .startofpacket
		.out_endofpacket   (st_bytes_to_packets_0_out_packets_stream_endofpacket),   //                   .endofpacket
		.in_ready          (sc_fifo_0_out_ready),                                    //    in_bytes_stream.ready
		.in_valid          (sc_fifo_0_out_valid),                                    //                   .valid
		.in_data           (sc_fifo_0_out_data)                                      //                   .data
	);

	altera_avalon_st_packets_to_bytes #(
		.CHANNEL_WIDTH (8),
		.ENCODING      (0)
	) st_packets_to_bytes_0 (
		.clk              (clk_clk),                                      //               clk.clk
		.reset_n          (reset_reset_n),                                //         clk_reset.reset_n
		.in_ready         (avalon_st_adapter_001_out_0_ready),            // in_packets_stream.ready
		.in_valid         (avalon_st_adapter_001_out_0_valid),            //                  .valid
		.in_data          (avalon_st_adapter_001_out_0_data),             //                  .data
		.in_channel       (avalon_st_adapter_001_out_0_channel),          //                  .channel
		.in_startofpacket (avalon_st_adapter_001_out_0_startofpacket),    //                  .startofpacket
		.in_endofpacket   (avalon_st_adapter_001_out_0_endofpacket),      //                  .endofpacket
		.out_ready        (st_packets_to_bytes_0_out_bytes_stream_ready), //  out_bytes_stream.ready
		.out_valid        (st_packets_to_bytes_0_out_bytes_stream_valid), //                  .valid
		.out_data         (st_packets_to_bytes_0_out_bytes_stream_data)   //                  .data
	);

	uart_to_bytes #(
		.CLOCK_FREQUENCY (100000000),
		.UART_BAUDRATE   (230400),
		.UART_STOPBIT    (1)
	) uart_to_bytes_0 (
		.clk       (clk_clk),                                      //  clock.clk
		.reset     (~reset_reset_n),                               //  reset.reset
		.txd       (uart_txd),                                     //   uart.txd
		.rxd       (uart_rxd),                                     //       .rxd
		.cts       (uart_cts),                                     //       .cts
		.rts       (uart_rts),                                     //       .rts
		.in_data   (st_packets_to_bytes_0_out_bytes_stream_data),  //   sink.data
		.in_ready  (st_packets_to_bytes_0_out_bytes_stream_ready), //       .ready
		.in_valid  (st_packets_to_bytes_0_out_bytes_stream_valid), //       .valid
		.out_data  (uart_to_bytes_0_source_data),                  // source.data
		.out_ready (uart_to_bytes_0_source_ready),                 //       .ready
		.out_valid (uart_to_bytes_0_source_valid)                  //       .valid
	);

	c4e_dvp_core_uart_to_avmm_bridge_avalon_st_adapter #(
		.inBitsPerSymbol (8),
		.inUsePackets    (1),
		.inDataWidth     (8),
		.inChannelWidth  (8),
		.inErrorWidth    (0),
		.inUseEmptyPort  (0),
		.inUseValid      (1),
		.inUseReady      (1),
		.inReadyLatency  (0),
		.outDataWidth    (8),
		.outChannelWidth (0),
		.outErrorWidth   (0),
		.outUseEmptyPort (0),
		.outUseValid     (1),
		.outUseReady     (1),
		.outReadyLatency (0)
	) avalon_st_adapter (
		.in_clk_0_clk        (clk_clk),                                                // in_clk_0.clk
		.in_rst_0_reset      (~reset_reset_n),                                         // in_rst_0.reset
		.in_0_data           (st_bytes_to_packets_0_out_packets_stream_data),          //     in_0.data
		.in_0_valid          (st_bytes_to_packets_0_out_packets_stream_valid),         //         .valid
		.in_0_ready          (st_bytes_to_packets_0_out_packets_stream_ready),         //         .ready
		.in_0_startofpacket  (st_bytes_to_packets_0_out_packets_stream_startofpacket), //         .startofpacket
		.in_0_endofpacket    (st_bytes_to_packets_0_out_packets_stream_endofpacket),   //         .endofpacket
		.in_0_channel        (st_bytes_to_packets_0_out_packets_stream_channel),       //         .channel
		.out_0_data          (avalon_st_adapter_out_0_data),                           //    out_0.data
		.out_0_valid         (avalon_st_adapter_out_0_valid),                          //         .valid
		.out_0_ready         (avalon_st_adapter_out_0_ready),                          //         .ready
		.out_0_startofpacket (avalon_st_adapter_out_0_startofpacket),                  //         .startofpacket
		.out_0_endofpacket   (avalon_st_adapter_out_0_endofpacket)                     //         .endofpacket
	);

	c4e_dvp_core_uart_to_avmm_bridge_avalon_st_adapter_001 #(
		.inBitsPerSymbol (8),
		.inUsePackets    (1),
		.inDataWidth     (8),
		.inChannelWidth  (0),
		.inErrorWidth    (0),
		.inUseEmptyPort  (0),
		.inUseValid      (1),
		.inUseReady      (1),
		.inReadyLatency  (0),
		.outDataWidth    (8),
		.outChannelWidth (8),
		.outErrorWidth   (0),
		.outUseEmptyPort (0),
		.outUseValid     (1),
		.outUseReady     (1),
		.outReadyLatency (0)
	) avalon_st_adapter_001 (
		.in_clk_0_clk        (clk_clk),                                      // in_clk_0.clk
		.in_rst_0_reset      (~reset_reset_n),                               // in_rst_0.reset
		.in_0_data           (packets_to_master_0_out_stream_data),          //     in_0.data
		.in_0_valid          (packets_to_master_0_out_stream_valid),         //         .valid
		.in_0_ready          (packets_to_master_0_out_stream_ready),         //         .ready
		.in_0_startofpacket  (packets_to_master_0_out_stream_startofpacket), //         .startofpacket
		.in_0_endofpacket    (packets_to_master_0_out_stream_endofpacket),   //         .endofpacket
		.out_0_data          (avalon_st_adapter_001_out_0_data),             //    out_0.data
		.out_0_valid         (avalon_st_adapter_001_out_0_valid),            //         .valid
		.out_0_ready         (avalon_st_adapter_001_out_0_ready),            //         .ready
		.out_0_startofpacket (avalon_st_adapter_001_out_0_startofpacket),    //         .startofpacket
		.out_0_endofpacket   (avalon_st_adapter_001_out_0_endofpacket),      //         .endofpacket
		.out_0_channel       (avalon_st_adapter_001_out_0_channel)           //         .channel
	);

endmodule
