// c4e_dvp_core.v

// Generated using ACDS version 20.1 720

`timescale 1 ps / 1 ps
module c4e_dvp_core (
		input  wire        clk_100m_clk,  // clk_100m.clk
		input  wire        clk_25m_clk,   //  clk_25m.clk
		input  wire        dvp_pclk,      //      dvp.pclk
		input  wire [7:0]  dvp_data,      //         .data
		input  wire        dvp_href,      //         .href
		input  wire        dvp_vsync,     //         .vsync
		output wire        dvp_reseto_n,  //         .reseto_n
		output wire        host_txd,      //     host.txd
		input  wire        host_rxd,      //         .rxd
		input  wire        host_cts,      //         .cts
		output wire        host_rts,      //         .rts
		output wire [3:0]  led_export,    //      led.export
		input  wire        reset_reset_n, //    reset.reset_n
		inout  wire        sccb_sck,      //     sccb.sck
		inout  wire        sccb_data,     //         .data
		output wire [12:0] sdr_addr,      //      sdr.addr
		output wire [1:0]  sdr_ba,        //         .ba
		output wire        sdr_cas_n,     //         .cas_n
		output wire        sdr_cke,       //         .cke
		output wire        sdr_cs_n,      //         .cs_n
		inout  wire [15:0] sdr_dq,        //         .dq
		output wire [1:0]  sdr_dqm,       //         .dqm
		output wire        sdr_ras_n,     //         .ras_n
		output wire        sdr_we_n,      //         .we_n
		input  wire        tmds_videoclk, //     tmds.videoclk
		input  wire        tmds_txclk,    //         .txclk
		output wire [2:0]  tmds_data,     //         .data
		output wire [2:0]  tmds_data_n,   //         .data_n
		output wire        tmds_clock,    //         .clock
		output wire        tmds_clock_n   //         .clock_n
	);

	wire  [31:0] uart_to_avmm_bridge_avm_readdata;                     // mm_interconnect_0:uart_to_avmm_bridge_avm_readdata -> uart_to_avmm_bridge:avm_readdata
	wire         uart_to_avmm_bridge_avm_waitrequest;                  // mm_interconnect_0:uart_to_avmm_bridge_avm_waitrequest -> uart_to_avmm_bridge:avm_waitrequest
	wire  [31:0] uart_to_avmm_bridge_avm_address;                      // uart_to_avmm_bridge:avm_address -> mm_interconnect_0:uart_to_avmm_bridge_avm_address
	wire         uart_to_avmm_bridge_avm_read;                         // uart_to_avmm_bridge:avm_read -> mm_interconnect_0:uart_to_avmm_bridge_avm_read
	wire   [3:0] uart_to_avmm_bridge_avm_byteenable;                   // uart_to_avmm_bridge:avm_byteenable -> mm_interconnect_0:uart_to_avmm_bridge_avm_byteenable
	wire         uart_to_avmm_bridge_avm_readdatavalid;                // mm_interconnect_0:uart_to_avmm_bridge_avm_readdatavalid -> uart_to_avmm_bridge:avm_readdatavalid
	wire         uart_to_avmm_bridge_avm_write;                        // uart_to_avmm_bridge:avm_write -> mm_interconnect_0:uart_to_avmm_bridge_avm_write
	wire  [31:0] uart_to_avmm_bridge_avm_writedata;                    // uart_to_avmm_bridge:avm_writedata -> mm_interconnect_0:uart_to_avmm_bridge_avm_writedata
	wire         vga_m1_waitrequest;                                   // mm_interconnect_0:vga_m1_waitrequest -> vga:avm_m1_waitrequest
	wire  [31:0] vga_m1_readdata;                                      // mm_interconnect_0:vga_m1_readdata -> vga:avm_m1_readdata
	wire  [31:0] vga_m1_address;                                       // vga:avm_m1_address -> mm_interconnect_0:vga_m1_address
	wire         vga_m1_read;                                          // vga:avm_m1_read -> mm_interconnect_0:vga_m1_read
	wire         vga_m1_readdatavalid;                                 // mm_interconnect_0:vga_m1_readdatavalid -> vga:avm_m1_readdatavalid
	wire   [8:0] vga_m1_burstcount;                                    // vga:avm_m1_burstcount -> mm_interconnect_0:vga_m1_burstcount
	wire         cam_m1_waitrequest;                                   // mm_interconnect_0:cam_m1_waitrequest -> cam:avm_m1_waitrequest
	wire  [31:0] cam_m1_address;                                       // cam:avm_m1_address -> mm_interconnect_0:cam_m1_address
	wire   [3:0] cam_m1_byteenable;                                    // cam:avm_m1_byteenable -> mm_interconnect_0:cam_m1_byteenable
	wire         cam_m1_write;                                         // cam:avm_m1_write -> mm_interconnect_0:cam_m1_write
	wire  [31:0] cam_m1_writedata;                                     // cam:avm_m1_writedata -> mm_interconnect_0:cam_m1_writedata
	wire   [8:0] cam_m1_burstcount;                                    // cam:avm_m1_burstcount -> mm_interconnect_0:cam_m1_burstcount
	wire  [31:0] mm_interconnect_0_peripheral_bridge_s0_readdata;      // peripheral_bridge:s0_readdata -> mm_interconnect_0:peripheral_bridge_s0_readdata
	wire         mm_interconnect_0_peripheral_bridge_s0_waitrequest;   // peripheral_bridge:s0_waitrequest -> mm_interconnect_0:peripheral_bridge_s0_waitrequest
	wire         mm_interconnect_0_peripheral_bridge_s0_debugaccess;   // mm_interconnect_0:peripheral_bridge_s0_debugaccess -> peripheral_bridge:s0_debugaccess
	wire   [9:0] mm_interconnect_0_peripheral_bridge_s0_address;       // mm_interconnect_0:peripheral_bridge_s0_address -> peripheral_bridge:s0_address
	wire         mm_interconnect_0_peripheral_bridge_s0_read;          // mm_interconnect_0:peripheral_bridge_s0_read -> peripheral_bridge:s0_read
	wire   [3:0] mm_interconnect_0_peripheral_bridge_s0_byteenable;    // mm_interconnect_0:peripheral_bridge_s0_byteenable -> peripheral_bridge:s0_byteenable
	wire         mm_interconnect_0_peripheral_bridge_s0_readdatavalid; // peripheral_bridge:s0_readdatavalid -> mm_interconnect_0:peripheral_bridge_s0_readdatavalid
	wire         mm_interconnect_0_peripheral_bridge_s0_write;         // mm_interconnect_0:peripheral_bridge_s0_write -> peripheral_bridge:s0_write
	wire  [31:0] mm_interconnect_0_peripheral_bridge_s0_writedata;     // mm_interconnect_0:peripheral_bridge_s0_writedata -> peripheral_bridge:s0_writedata
	wire   [0:0] mm_interconnect_0_peripheral_bridge_s0_burstcount;    // mm_interconnect_0:peripheral_bridge_s0_burstcount -> peripheral_bridge:s0_burstcount
	wire         mm_interconnect_0_sdram_s1_chipselect;                // mm_interconnect_0:sdram_s1_chipselect -> sdram:az_cs
	wire  [15:0] mm_interconnect_0_sdram_s1_readdata;                  // sdram:za_data -> mm_interconnect_0:sdram_s1_readdata
	wire         mm_interconnect_0_sdram_s1_waitrequest;               // sdram:za_waitrequest -> mm_interconnect_0:sdram_s1_waitrequest
	wire  [23:0] mm_interconnect_0_sdram_s1_address;                   // mm_interconnect_0:sdram_s1_address -> sdram:az_addr
	wire         mm_interconnect_0_sdram_s1_read;                      // mm_interconnect_0:sdram_s1_read -> sdram:az_rd_n
	wire   [1:0] mm_interconnect_0_sdram_s1_byteenable;                // mm_interconnect_0:sdram_s1_byteenable -> sdram:az_be_n
	wire         mm_interconnect_0_sdram_s1_readdatavalid;             // sdram:za_valid -> mm_interconnect_0:sdram_s1_readdatavalid
	wire         mm_interconnect_0_sdram_s1_write;                     // mm_interconnect_0:sdram_s1_write -> sdram:az_wr_n
	wire  [15:0] mm_interconnect_0_sdram_s1_writedata;                 // mm_interconnect_0:sdram_s1_writedata -> sdram:az_data
	wire         peripheral_bridge_m0_waitrequest;                     // mm_interconnect_1:peripheral_bridge_m0_waitrequest -> peripheral_bridge:m0_waitrequest
	wire  [31:0] peripheral_bridge_m0_readdata;                        // mm_interconnect_1:peripheral_bridge_m0_readdata -> peripheral_bridge:m0_readdata
	wire         peripheral_bridge_m0_debugaccess;                     // peripheral_bridge:m0_debugaccess -> mm_interconnect_1:peripheral_bridge_m0_debugaccess
	wire   [9:0] peripheral_bridge_m0_address;                         // peripheral_bridge:m0_address -> mm_interconnect_1:peripheral_bridge_m0_address
	wire         peripheral_bridge_m0_read;                            // peripheral_bridge:m0_read -> mm_interconnect_1:peripheral_bridge_m0_read
	wire   [3:0] peripheral_bridge_m0_byteenable;                      // peripheral_bridge:m0_byteenable -> mm_interconnect_1:peripheral_bridge_m0_byteenable
	wire         peripheral_bridge_m0_readdatavalid;                   // mm_interconnect_1:peripheral_bridge_m0_readdatavalid -> peripheral_bridge:m0_readdatavalid
	wire  [31:0] peripheral_bridge_m0_writedata;                       // peripheral_bridge:m0_writedata -> mm_interconnect_1:peripheral_bridge_m0_writedata
	wire         peripheral_bridge_m0_write;                           // peripheral_bridge:m0_write -> mm_interconnect_1:peripheral_bridge_m0_write
	wire   [0:0] peripheral_bridge_m0_burstcount;                      // peripheral_bridge:m0_burstcount -> mm_interconnect_1:peripheral_bridge_m0_burstcount
	wire  [31:0] mm_interconnect_1_sysid_control_slave_readdata;       // sysid:readdata -> mm_interconnect_1:sysid_control_slave_readdata
	wire   [0:0] mm_interconnect_1_sysid_control_slave_address;        // mm_interconnect_1:sysid_control_slave_address -> sysid:address
	wire  [31:0] mm_interconnect_1_vga_csr_readdata;                   // vga:avs_csr_readdata -> mm_interconnect_1:vga_csr_readdata
	wire   [1:0] mm_interconnect_1_vga_csr_address;                    // mm_interconnect_1:vga_csr_address -> vga:avs_csr_address
	wire         mm_interconnect_1_vga_csr_read;                       // mm_interconnect_1:vga_csr_read -> vga:avs_csr_read
	wire         mm_interconnect_1_vga_csr_write;                      // mm_interconnect_1:vga_csr_write -> vga:avs_csr_write
	wire  [31:0] mm_interconnect_1_vga_csr_writedata;                  // mm_interconnect_1:vga_csr_writedata -> vga:avs_csr_writedata
	wire         mm_interconnect_1_led_s1_chipselect;                  // mm_interconnect_1:led_s1_chipselect -> led:chipselect
	wire  [31:0] mm_interconnect_1_led_s1_readdata;                    // led:readdata -> mm_interconnect_1:led_s1_readdata
	wire   [1:0] mm_interconnect_1_led_s1_address;                     // mm_interconnect_1:led_s1_address -> led:address
	wire         mm_interconnect_1_led_s1_write;                       // mm_interconnect_1:led_s1_write -> led:write_n
	wire  [31:0] mm_interconnect_1_led_s1_writedata;                   // mm_interconnect_1:led_s1_writedata -> led:writedata
	wire  [31:0] mm_interconnect_1_cam_s1_readdata;                    // cam:avs_s1_readdata -> mm_interconnect_1:cam_s1_readdata
	wire         mm_interconnect_1_cam_s1_waitrequest;                 // cam:avs_s1_waitrequest -> mm_interconnect_1:cam_s1_waitrequest
	wire   [1:0] mm_interconnect_1_cam_s1_address;                     // mm_interconnect_1:cam_s1_address -> cam:avs_s1_address
	wire         mm_interconnect_1_cam_s1_read;                        // mm_interconnect_1:cam_s1_read -> cam:avs_s1_read
	wire         mm_interconnect_1_cam_s1_write;                       // mm_interconnect_1:cam_s1_write -> cam:avs_s1_write
	wire  [31:0] mm_interconnect_1_cam_s1_writedata;                   // mm_interconnect_1:cam_s1_writedata -> cam:avs_s1_writedata
	wire         rst_controller_reset_out_reset;                       // rst_controller:reset_out -> [cam:csi_global_reset, led:reset_n, mm_interconnect_0:peripheral_bridge_reset_reset_bridge_in_reset_reset, mm_interconnect_1:peripheral_bridge_reset_reset_bridge_in_reset_reset, peripheral_bridge:reset, sysid:reset_n, vga:csi_csr_reset]
	wire         rst_controller_001_reset_out_reset;                   // rst_controller_001:reset_out -> [mm_interconnect_0:uart_to_avmm_bridge_reset_reset_bridge_in_reset_reset, sdram:reset_n, uart_to_avmm_bridge:reset_reset_n]
	wire         rst_controller_002_reset_out_reset;                   // rst_controller_002:reset_out -> mm_interconnect_0:vga_reset_reset_bridge_in_reset_reset

	peridot_cam #(
		.AVM_CLOCKFREQ     (100000000),
		.AVS_CLOCKFREQ     (25000000),
		.BURSTCOUNT_WIDTH  (8),
		.TRANSCYCLE_WIDTH  (22),
		.DVP_FIFO_DEPTH    (12),
		.DVP_BYTESWAP      ("OFF"),
		.USE_SCCBINTERFACE ("ON"),
		.USE_PERIDOT_I2C   ("OFF"),
		.SCCB_CLOCKFREQ    (400000)
	) cam (
		.csi_global_clk     (clk_25m_clk),                          // s1_clock.clk
		.csi_global_reset   (rst_controller_reset_out_reset),       // s1_reset.reset
		.avs_s1_address     (mm_interconnect_1_cam_s1_address),     //       s1.address
		.avs_s1_write       (mm_interconnect_1_cam_s1_write),       //         .write
		.avs_s1_writedata   (mm_interconnect_1_cam_s1_writedata),   //         .writedata
		.avs_s1_read        (mm_interconnect_1_cam_s1_read),        //         .read
		.avs_s1_readdata    (mm_interconnect_1_cam_s1_readdata),    //         .readdata
		.avs_s1_waitrequest (mm_interconnect_1_cam_s1_waitrequest), //         .waitrequest
		.avs_s1_irq         (),                                     //   irq_s1.irq
		.avm_m1_clk         (clk_100m_clk),                         // m1_clock.clk
		.avm_m1_address     (cam_m1_address),                       //       m1.address
		.avm_m1_write       (cam_m1_write),                         //         .write
		.avm_m1_writedata   (cam_m1_writedata),                     //         .writedata
		.avm_m1_byteenable  (cam_m1_byteenable),                    //         .byteenable
		.avm_m1_waitrequest (cam_m1_waitrequest),                   //         .waitrequest
		.avm_m1_burstcount  (cam_m1_burstcount),                    //         .burstcount
		.cam_clk            (dvp_pclk),                             //      dvp.pclk
		.cam_data           (dvp_data),                             //         .data
		.cam_href           (dvp_href),                             //         .href
		.cam_vsync          (dvp_vsync),                            //         .vsync
		.cam_reset_n        (dvp_reseto_n),                         //         .reseto_n
		.sccb_sck           (sccb_sck),                             //     sccb.sck
		.sccb_data          (sccb_data)                             //         .data
	);

	c4e_dvp_core_led led (
		.clk        (clk_25m_clk),                         //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),     //               reset.reset_n
		.address    (mm_interconnect_1_led_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_1_led_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_1_led_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_1_led_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_1_led_s1_readdata),   //                    .readdata
		.out_port   (led_export)                           // external_connection.export
	);

	altera_avalon_mm_bridge #(
		.DATA_WIDTH        (32),
		.SYMBOL_WIDTH      (8),
		.HDL_ADDR_WIDTH    (10),
		.BURSTCOUNT_WIDTH  (1),
		.PIPELINE_COMMAND  (1),
		.PIPELINE_RESPONSE (1)
	) peripheral_bridge (
		.clk              (clk_25m_clk),                                          //   clk.clk
		.reset            (rst_controller_reset_out_reset),                       // reset.reset
		.s0_waitrequest   (mm_interconnect_0_peripheral_bridge_s0_waitrequest),   //    s0.waitrequest
		.s0_readdata      (mm_interconnect_0_peripheral_bridge_s0_readdata),      //      .readdata
		.s0_readdatavalid (mm_interconnect_0_peripheral_bridge_s0_readdatavalid), //      .readdatavalid
		.s0_burstcount    (mm_interconnect_0_peripheral_bridge_s0_burstcount),    //      .burstcount
		.s0_writedata     (mm_interconnect_0_peripheral_bridge_s0_writedata),     //      .writedata
		.s0_address       (mm_interconnect_0_peripheral_bridge_s0_address),       //      .address
		.s0_write         (mm_interconnect_0_peripheral_bridge_s0_write),         //      .write
		.s0_read          (mm_interconnect_0_peripheral_bridge_s0_read),          //      .read
		.s0_byteenable    (mm_interconnect_0_peripheral_bridge_s0_byteenable),    //      .byteenable
		.s0_debugaccess   (mm_interconnect_0_peripheral_bridge_s0_debugaccess),   //      .debugaccess
		.m0_waitrequest   (peripheral_bridge_m0_waitrequest),                     //    m0.waitrequest
		.m0_readdata      (peripheral_bridge_m0_readdata),                        //      .readdata
		.m0_readdatavalid (peripheral_bridge_m0_readdatavalid),                   //      .readdatavalid
		.m0_burstcount    (peripheral_bridge_m0_burstcount),                      //      .burstcount
		.m0_writedata     (peripheral_bridge_m0_writedata),                       //      .writedata
		.m0_address       (peripheral_bridge_m0_address),                         //      .address
		.m0_write         (peripheral_bridge_m0_write),                           //      .write
		.m0_read          (peripheral_bridge_m0_read),                            //      .read
		.m0_byteenable    (peripheral_bridge_m0_byteenable),                      //      .byteenable
		.m0_debugaccess   (peripheral_bridge_m0_debugaccess),                     //      .debugaccess
		.s0_response      (),                                                     // (terminated)
		.m0_response      (2'b00)                                                 // (terminated)
	);

	c4e_dvp_core_sdram sdram (
		.clk            (clk_100m_clk),                             //   clk.clk
		.reset_n        (~rst_controller_001_reset_out_reset),      // reset.reset_n
		.az_addr        (mm_interconnect_0_sdram_s1_address),       //    s1.address
		.az_be_n        (~mm_interconnect_0_sdram_s1_byteenable),   //      .byteenable_n
		.az_cs          (mm_interconnect_0_sdram_s1_chipselect),    //      .chipselect
		.az_data        (mm_interconnect_0_sdram_s1_writedata),     //      .writedata
		.az_rd_n        (~mm_interconnect_0_sdram_s1_read),         //      .read_n
		.az_wr_n        (~mm_interconnect_0_sdram_s1_write),        //      .write_n
		.za_data        (mm_interconnect_0_sdram_s1_readdata),      //      .readdata
		.za_valid       (mm_interconnect_0_sdram_s1_readdatavalid), //      .readdatavalid
		.za_waitrequest (mm_interconnect_0_sdram_s1_waitrequest),   //      .waitrequest
		.zs_addr        (sdr_addr),                                 //  wire.export
		.zs_ba          (sdr_ba),                                   //      .export
		.zs_cas_n       (sdr_cas_n),                                //      .export
		.zs_cke         (sdr_cke),                                  //      .export
		.zs_cs_n        (sdr_cs_n),                                 //      .export
		.zs_dq          (sdr_dq),                                   //      .export
		.zs_dqm         (sdr_dqm),                                  //      .export
		.zs_ras_n       (sdr_ras_n),                                //      .export
		.zs_we_n        (sdr_we_n)                                  //      .export
	);

	c4e_dvp_core_sysid sysid (
		.clock    (clk_25m_clk),                                    //           clk.clk
		.reset_n  (~rst_controller_reset_out_reset),                //         reset.reset_n
		.readdata (mm_interconnect_1_sysid_control_slave_readdata), // control_slave.readdata
		.address  (mm_interconnect_1_sysid_control_slave_address)   //              .address
	);

	c4e_dvp_core_uart_to_avmm_bridge uart_to_avmm_bridge (
		.avm_address       (uart_to_avmm_bridge_avm_address),       //   avm.address
		.avm_readdata      (uart_to_avmm_bridge_avm_readdata),      //      .readdata
		.avm_read          (uart_to_avmm_bridge_avm_read),          //      .read
		.avm_write         (uart_to_avmm_bridge_avm_write),         //      .write
		.avm_writedata     (uart_to_avmm_bridge_avm_writedata),     //      .writedata
		.avm_waitrequest   (uart_to_avmm_bridge_avm_waitrequest),   //      .waitrequest
		.avm_readdatavalid (uart_to_avmm_bridge_avm_readdatavalid), //      .readdatavalid
		.avm_byteenable    (uart_to_avmm_bridge_avm_byteenable),    //      .byteenable
		.clk_clk           (clk_100m_clk),                          //   clk.clk
		.reset_reset_n     (~rst_controller_001_reset_out_reset),   // reset.reset_n
		.uart_txd          (host_txd),                              //  uart.txd
		.uart_rxd          (host_rxd),                              //      .rxd
		.uart_cts          (host_cts),                              //      .cts
		.uart_rts          (host_rts)                               //      .rts
	);

	peridot_vga #(
		.DEVICE_FAMILY       ("Cyclone IV E"),
		.FIFORESETCOUNT      (10),
		.FIFODEPTH_WIDTH     (10),
		.VIDEO_INTERFACE     ("DVI"),
		.VGACLOCK_FREQUENCY  (65000000),
		.H_TOTAL             (1344),
		.H_SYNC              (136),
		.H_BACKP             (160),
		.H_ACTIVE            (1024),
		.V_TOTAL             (806),
		.V_SYNC              (6),
		.V_BACKP             (29),
		.V_ACTIVE            (768),
		.USE_AUDIOSTREAM     ("OFF"),
		.BURSTCOUNT_WIDTH    (8),
		.LINEOFFSETBYTES     (2560),
		.PIXEL_DATAORDER     ("BYTE"),
		.PIXEL_COLORORDER    ("YUV422"),
		.PCMSAMPLE_FREQUENCY (44100)
	) vga (
		.csi_csr_clk          (clk_25m_clk),                         // csr_clk.clk
		.csi_csr_reset        (rst_controller_reset_out_reset),      //   reset.reset
		.avs_csr_address      (mm_interconnect_1_vga_csr_address),   //     csr.address
		.avs_csr_read         (mm_interconnect_1_vga_csr_read),      //        .read
		.avs_csr_readdata     (mm_interconnect_1_vga_csr_readdata),  //        .readdata
		.avs_csr_write        (mm_interconnect_1_vga_csr_write),     //        .write
		.avs_csr_writedata    (mm_interconnect_1_vga_csr_writedata), //        .writedata
		.ins_csr_irq          (),                                    // irq_csr.irq
		.csi_m1_clk           (clk_100m_clk),                        //  m1_clk.clk
		.avm_m1_waitrequest   (vga_m1_waitrequest),                  //      m1.waitrequest
		.avm_m1_address       (vga_m1_address),                      //        .address
		.avm_m1_read          (vga_m1_read),                         //        .read
		.avm_m1_readdata      (vga_m1_readdata),                     //        .readdata
		.avm_m1_readdatavalid (vga_m1_readdatavalid),                //        .readdatavalid
		.avm_m1_burstcount    (vga_m1_burstcount),                   //        .burstcount
		.coe_ser_clk          (tmds_videoclk),                       //    tmds.videoclk
		.coe_ser_x5clk        (tmds_txclk),                          //        .txclk
		.coe_ser_data         (tmds_data),                           //        .data
		.coe_ser_data_n       (tmds_data_n),                         //        .data_n
		.coe_ser_clock        (tmds_clock),                          //        .clock
		.coe_ser_clock_n      (tmds_clock_n),                        //        .clock_n
		.coe_pcm_fs           (1'b0),                                // (terminated)
		.coe_pcm_l            (24'b000000000000000000000000),        // (terminated)
		.coe_pcm_r            (24'b000000000000000000000000),        // (terminated)
		.coe_vga_clk          (1'b0),                                // (terminated)
		.coe_vga_active       (),                                    // (terminated)
		.coe_vga_rout         (),                                    // (terminated)
		.coe_vga_gout         (),                                    // (terminated)
		.coe_vga_bout         (),                                    // (terminated)
		.coe_vga_hsync_n      (),                                    // (terminated)
		.coe_vga_vsync_n      (),                                    // (terminated)
		.coe_vga_csync_n      ()                                     // (terminated)
	);

	c4e_dvp_core_mm_interconnect_0 mm_interconnect_0 (
		.core_clk_clk_clk                                      (clk_100m_clk),                                         //                                    core_clk_clk.clk
		.peri_clk_clk_clk                                      (clk_25m_clk),                                          //                                    peri_clk_clk.clk
		.peripheral_bridge_reset_reset_bridge_in_reset_reset   (rst_controller_reset_out_reset),                       //   peripheral_bridge_reset_reset_bridge_in_reset.reset
		.uart_to_avmm_bridge_reset_reset_bridge_in_reset_reset (rst_controller_001_reset_out_reset),                   // uart_to_avmm_bridge_reset_reset_bridge_in_reset.reset
		.vga_reset_reset_bridge_in_reset_reset                 (rst_controller_002_reset_out_reset),                   //                 vga_reset_reset_bridge_in_reset.reset
		.cam_m1_address                                        (cam_m1_address),                                       //                                          cam_m1.address
		.cam_m1_waitrequest                                    (cam_m1_waitrequest),                                   //                                                .waitrequest
		.cam_m1_burstcount                                     (cam_m1_burstcount),                                    //                                                .burstcount
		.cam_m1_byteenable                                     (cam_m1_byteenable),                                    //                                                .byteenable
		.cam_m1_write                                          (cam_m1_write),                                         //                                                .write
		.cam_m1_writedata                                      (cam_m1_writedata),                                     //                                                .writedata
		.uart_to_avmm_bridge_avm_address                       (uart_to_avmm_bridge_avm_address),                      //                         uart_to_avmm_bridge_avm.address
		.uart_to_avmm_bridge_avm_waitrequest                   (uart_to_avmm_bridge_avm_waitrequest),                  //                                                .waitrequest
		.uart_to_avmm_bridge_avm_byteenable                    (uart_to_avmm_bridge_avm_byteenable),                   //                                                .byteenable
		.uart_to_avmm_bridge_avm_read                          (uart_to_avmm_bridge_avm_read),                         //                                                .read
		.uart_to_avmm_bridge_avm_readdata                      (uart_to_avmm_bridge_avm_readdata),                     //                                                .readdata
		.uart_to_avmm_bridge_avm_readdatavalid                 (uart_to_avmm_bridge_avm_readdatavalid),                //                                                .readdatavalid
		.uart_to_avmm_bridge_avm_write                         (uart_to_avmm_bridge_avm_write),                        //                                                .write
		.uart_to_avmm_bridge_avm_writedata                     (uart_to_avmm_bridge_avm_writedata),                    //                                                .writedata
		.vga_m1_address                                        (vga_m1_address),                                       //                                          vga_m1.address
		.vga_m1_waitrequest                                    (vga_m1_waitrequest),                                   //                                                .waitrequest
		.vga_m1_burstcount                                     (vga_m1_burstcount),                                    //                                                .burstcount
		.vga_m1_read                                           (vga_m1_read),                                          //                                                .read
		.vga_m1_readdata                                       (vga_m1_readdata),                                      //                                                .readdata
		.vga_m1_readdatavalid                                  (vga_m1_readdatavalid),                                 //                                                .readdatavalid
		.peripheral_bridge_s0_address                          (mm_interconnect_0_peripheral_bridge_s0_address),       //                            peripheral_bridge_s0.address
		.peripheral_bridge_s0_write                            (mm_interconnect_0_peripheral_bridge_s0_write),         //                                                .write
		.peripheral_bridge_s0_read                             (mm_interconnect_0_peripheral_bridge_s0_read),          //                                                .read
		.peripheral_bridge_s0_readdata                         (mm_interconnect_0_peripheral_bridge_s0_readdata),      //                                                .readdata
		.peripheral_bridge_s0_writedata                        (mm_interconnect_0_peripheral_bridge_s0_writedata),     //                                                .writedata
		.peripheral_bridge_s0_burstcount                       (mm_interconnect_0_peripheral_bridge_s0_burstcount),    //                                                .burstcount
		.peripheral_bridge_s0_byteenable                       (mm_interconnect_0_peripheral_bridge_s0_byteenable),    //                                                .byteenable
		.peripheral_bridge_s0_readdatavalid                    (mm_interconnect_0_peripheral_bridge_s0_readdatavalid), //                                                .readdatavalid
		.peripheral_bridge_s0_waitrequest                      (mm_interconnect_0_peripheral_bridge_s0_waitrequest),   //                                                .waitrequest
		.peripheral_bridge_s0_debugaccess                      (mm_interconnect_0_peripheral_bridge_s0_debugaccess),   //                                                .debugaccess
		.sdram_s1_address                                      (mm_interconnect_0_sdram_s1_address),                   //                                        sdram_s1.address
		.sdram_s1_write                                        (mm_interconnect_0_sdram_s1_write),                     //                                                .write
		.sdram_s1_read                                         (mm_interconnect_0_sdram_s1_read),                      //                                                .read
		.sdram_s1_readdata                                     (mm_interconnect_0_sdram_s1_readdata),                  //                                                .readdata
		.sdram_s1_writedata                                    (mm_interconnect_0_sdram_s1_writedata),                 //                                                .writedata
		.sdram_s1_byteenable                                   (mm_interconnect_0_sdram_s1_byteenable),                //                                                .byteenable
		.sdram_s1_readdatavalid                                (mm_interconnect_0_sdram_s1_readdatavalid),             //                                                .readdatavalid
		.sdram_s1_waitrequest                                  (mm_interconnect_0_sdram_s1_waitrequest),               //                                                .waitrequest
		.sdram_s1_chipselect                                   (mm_interconnect_0_sdram_s1_chipselect)                 //                                                .chipselect
	);

	c4e_dvp_core_mm_interconnect_1 mm_interconnect_1 (
		.peri_clk_clk_clk                                    (clk_25m_clk),                                    //                                  peri_clk_clk.clk
		.peripheral_bridge_reset_reset_bridge_in_reset_reset (rst_controller_reset_out_reset),                 // peripheral_bridge_reset_reset_bridge_in_reset.reset
		.peripheral_bridge_m0_address                        (peripheral_bridge_m0_address),                   //                          peripheral_bridge_m0.address
		.peripheral_bridge_m0_waitrequest                    (peripheral_bridge_m0_waitrequest),               //                                              .waitrequest
		.peripheral_bridge_m0_burstcount                     (peripheral_bridge_m0_burstcount),                //                                              .burstcount
		.peripheral_bridge_m0_byteenable                     (peripheral_bridge_m0_byteenable),                //                                              .byteenable
		.peripheral_bridge_m0_read                           (peripheral_bridge_m0_read),                      //                                              .read
		.peripheral_bridge_m0_readdata                       (peripheral_bridge_m0_readdata),                  //                                              .readdata
		.peripheral_bridge_m0_readdatavalid                  (peripheral_bridge_m0_readdatavalid),             //                                              .readdatavalid
		.peripheral_bridge_m0_write                          (peripheral_bridge_m0_write),                     //                                              .write
		.peripheral_bridge_m0_writedata                      (peripheral_bridge_m0_writedata),                 //                                              .writedata
		.peripheral_bridge_m0_debugaccess                    (peripheral_bridge_m0_debugaccess),               //                                              .debugaccess
		.cam_s1_address                                      (mm_interconnect_1_cam_s1_address),               //                                        cam_s1.address
		.cam_s1_write                                        (mm_interconnect_1_cam_s1_write),                 //                                              .write
		.cam_s1_read                                         (mm_interconnect_1_cam_s1_read),                  //                                              .read
		.cam_s1_readdata                                     (mm_interconnect_1_cam_s1_readdata),              //                                              .readdata
		.cam_s1_writedata                                    (mm_interconnect_1_cam_s1_writedata),             //                                              .writedata
		.cam_s1_waitrequest                                  (mm_interconnect_1_cam_s1_waitrequest),           //                                              .waitrequest
		.led_s1_address                                      (mm_interconnect_1_led_s1_address),               //                                        led_s1.address
		.led_s1_write                                        (mm_interconnect_1_led_s1_write),                 //                                              .write
		.led_s1_readdata                                     (mm_interconnect_1_led_s1_readdata),              //                                              .readdata
		.led_s1_writedata                                    (mm_interconnect_1_led_s1_writedata),             //                                              .writedata
		.led_s1_chipselect                                   (mm_interconnect_1_led_s1_chipselect),            //                                              .chipselect
		.sysid_control_slave_address                         (mm_interconnect_1_sysid_control_slave_address),  //                           sysid_control_slave.address
		.sysid_control_slave_readdata                        (mm_interconnect_1_sysid_control_slave_readdata), //                                              .readdata
		.vga_csr_address                                     (mm_interconnect_1_vga_csr_address),              //                                       vga_csr.address
		.vga_csr_write                                       (mm_interconnect_1_vga_csr_write),                //                                              .write
		.vga_csr_read                                        (mm_interconnect_1_vga_csr_read),                 //                                              .read
		.vga_csr_readdata                                    (mm_interconnect_1_vga_csr_readdata),             //                                              .readdata
		.vga_csr_writedata                                   (mm_interconnect_1_vga_csr_writedata)             //                                              .writedata
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS          (1),
		.OUTPUT_RESET_SYNC_EDGES   ("deassert"),
		.SYNC_DEPTH                (2),
		.RESET_REQUEST_PRESENT     (0),
		.RESET_REQ_WAIT_TIME       (1),
		.MIN_RST_ASSERTION_TIME    (3),
		.RESET_REQ_EARLY_DSRT_TIME (1),
		.USE_RESET_REQUEST_IN0     (0),
		.USE_RESET_REQUEST_IN1     (0),
		.USE_RESET_REQUEST_IN2     (0),
		.USE_RESET_REQUEST_IN3     (0),
		.USE_RESET_REQUEST_IN4     (0),
		.USE_RESET_REQUEST_IN5     (0),
		.USE_RESET_REQUEST_IN6     (0),
		.USE_RESET_REQUEST_IN7     (0),
		.USE_RESET_REQUEST_IN8     (0),
		.USE_RESET_REQUEST_IN9     (0),
		.USE_RESET_REQUEST_IN10    (0),
		.USE_RESET_REQUEST_IN11    (0),
		.USE_RESET_REQUEST_IN12    (0),
		.USE_RESET_REQUEST_IN13    (0),
		.USE_RESET_REQUEST_IN14    (0),
		.USE_RESET_REQUEST_IN15    (0),
		.ADAPT_RESET_REQUEST       (0)
	) rst_controller (
		.reset_in0      (~reset_reset_n),                 // reset_in0.reset
		.clk            (clk_25m_clk),                    //       clk.clk
		.reset_out      (rst_controller_reset_out_reset), // reset_out.reset
		.reset_req      (),                               // (terminated)
		.reset_req_in0  (1'b0),                           // (terminated)
		.reset_in1      (1'b0),                           // (terminated)
		.reset_req_in1  (1'b0),                           // (terminated)
		.reset_in2      (1'b0),                           // (terminated)
		.reset_req_in2  (1'b0),                           // (terminated)
		.reset_in3      (1'b0),                           // (terminated)
		.reset_req_in3  (1'b0),                           // (terminated)
		.reset_in4      (1'b0),                           // (terminated)
		.reset_req_in4  (1'b0),                           // (terminated)
		.reset_in5      (1'b0),                           // (terminated)
		.reset_req_in5  (1'b0),                           // (terminated)
		.reset_in6      (1'b0),                           // (terminated)
		.reset_req_in6  (1'b0),                           // (terminated)
		.reset_in7      (1'b0),                           // (terminated)
		.reset_req_in7  (1'b0),                           // (terminated)
		.reset_in8      (1'b0),                           // (terminated)
		.reset_req_in8  (1'b0),                           // (terminated)
		.reset_in9      (1'b0),                           // (terminated)
		.reset_req_in9  (1'b0),                           // (terminated)
		.reset_in10     (1'b0),                           // (terminated)
		.reset_req_in10 (1'b0),                           // (terminated)
		.reset_in11     (1'b0),                           // (terminated)
		.reset_req_in11 (1'b0),                           // (terminated)
		.reset_in12     (1'b0),                           // (terminated)
		.reset_req_in12 (1'b0),                           // (terminated)
		.reset_in13     (1'b0),                           // (terminated)
		.reset_req_in13 (1'b0),                           // (terminated)
		.reset_in14     (1'b0),                           // (terminated)
		.reset_req_in14 (1'b0),                           // (terminated)
		.reset_in15     (1'b0),                           // (terminated)
		.reset_req_in15 (1'b0)                            // (terminated)
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS          (1),
		.OUTPUT_RESET_SYNC_EDGES   ("deassert"),
		.SYNC_DEPTH                (2),
		.RESET_REQUEST_PRESENT     (0),
		.RESET_REQ_WAIT_TIME       (1),
		.MIN_RST_ASSERTION_TIME    (3),
		.RESET_REQ_EARLY_DSRT_TIME (1),
		.USE_RESET_REQUEST_IN0     (0),
		.USE_RESET_REQUEST_IN1     (0),
		.USE_RESET_REQUEST_IN2     (0),
		.USE_RESET_REQUEST_IN3     (0),
		.USE_RESET_REQUEST_IN4     (0),
		.USE_RESET_REQUEST_IN5     (0),
		.USE_RESET_REQUEST_IN6     (0),
		.USE_RESET_REQUEST_IN7     (0),
		.USE_RESET_REQUEST_IN8     (0),
		.USE_RESET_REQUEST_IN9     (0),
		.USE_RESET_REQUEST_IN10    (0),
		.USE_RESET_REQUEST_IN11    (0),
		.USE_RESET_REQUEST_IN12    (0),
		.USE_RESET_REQUEST_IN13    (0),
		.USE_RESET_REQUEST_IN14    (0),
		.USE_RESET_REQUEST_IN15    (0),
		.ADAPT_RESET_REQUEST       (0)
	) rst_controller_001 (
		.reset_in0      (~reset_reset_n),                     // reset_in0.reset
		.clk            (clk_100m_clk),                       //       clk.clk
		.reset_out      (rst_controller_001_reset_out_reset), // reset_out.reset
		.reset_req      (),                                   // (terminated)
		.reset_req_in0  (1'b0),                               // (terminated)
		.reset_in1      (1'b0),                               // (terminated)
		.reset_req_in1  (1'b0),                               // (terminated)
		.reset_in2      (1'b0),                               // (terminated)
		.reset_req_in2  (1'b0),                               // (terminated)
		.reset_in3      (1'b0),                               // (terminated)
		.reset_req_in3  (1'b0),                               // (terminated)
		.reset_in4      (1'b0),                               // (terminated)
		.reset_req_in4  (1'b0),                               // (terminated)
		.reset_in5      (1'b0),                               // (terminated)
		.reset_req_in5  (1'b0),                               // (terminated)
		.reset_in6      (1'b0),                               // (terminated)
		.reset_req_in6  (1'b0),                               // (terminated)
		.reset_in7      (1'b0),                               // (terminated)
		.reset_req_in7  (1'b0),                               // (terminated)
		.reset_in8      (1'b0),                               // (terminated)
		.reset_req_in8  (1'b0),                               // (terminated)
		.reset_in9      (1'b0),                               // (terminated)
		.reset_req_in9  (1'b0),                               // (terminated)
		.reset_in10     (1'b0),                               // (terminated)
		.reset_req_in10 (1'b0),                               // (terminated)
		.reset_in11     (1'b0),                               // (terminated)
		.reset_req_in11 (1'b0),                               // (terminated)
		.reset_in12     (1'b0),                               // (terminated)
		.reset_req_in12 (1'b0),                               // (terminated)
		.reset_in13     (1'b0),                               // (terminated)
		.reset_req_in13 (1'b0),                               // (terminated)
		.reset_in14     (1'b0),                               // (terminated)
		.reset_req_in14 (1'b0),                               // (terminated)
		.reset_in15     (1'b0),                               // (terminated)
		.reset_req_in15 (1'b0)                                // (terminated)
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS          (1),
		.OUTPUT_RESET_SYNC_EDGES   ("deassert"),
		.SYNC_DEPTH                (2),
		.RESET_REQUEST_PRESENT     (0),
		.RESET_REQ_WAIT_TIME       (1),
		.MIN_RST_ASSERTION_TIME    (3),
		.RESET_REQ_EARLY_DSRT_TIME (1),
		.USE_RESET_REQUEST_IN0     (0),
		.USE_RESET_REQUEST_IN1     (0),
		.USE_RESET_REQUEST_IN2     (0),
		.USE_RESET_REQUEST_IN3     (0),
		.USE_RESET_REQUEST_IN4     (0),
		.USE_RESET_REQUEST_IN5     (0),
		.USE_RESET_REQUEST_IN6     (0),
		.USE_RESET_REQUEST_IN7     (0),
		.USE_RESET_REQUEST_IN8     (0),
		.USE_RESET_REQUEST_IN9     (0),
		.USE_RESET_REQUEST_IN10    (0),
		.USE_RESET_REQUEST_IN11    (0),
		.USE_RESET_REQUEST_IN12    (0),
		.USE_RESET_REQUEST_IN13    (0),
		.USE_RESET_REQUEST_IN14    (0),
		.USE_RESET_REQUEST_IN15    (0),
		.ADAPT_RESET_REQUEST       (0)
	) rst_controller_002 (
		.reset_in0      (~reset_reset_n),                     // reset_in0.reset
		.clk            (clk_100m_clk),                       //       clk.clk
		.reset_out      (rst_controller_002_reset_out_reset), // reset_out.reset
		.reset_req      (),                                   // (terminated)
		.reset_req_in0  (1'b0),                               // (terminated)
		.reset_in1      (1'b0),                               // (terminated)
		.reset_req_in1  (1'b0),                               // (terminated)
		.reset_in2      (1'b0),                               // (terminated)
		.reset_req_in2  (1'b0),                               // (terminated)
		.reset_in3      (1'b0),                               // (terminated)
		.reset_req_in3  (1'b0),                               // (terminated)
		.reset_in4      (1'b0),                               // (terminated)
		.reset_req_in4  (1'b0),                               // (terminated)
		.reset_in5      (1'b0),                               // (terminated)
		.reset_req_in5  (1'b0),                               // (terminated)
		.reset_in6      (1'b0),                               // (terminated)
		.reset_req_in6  (1'b0),                               // (terminated)
		.reset_in7      (1'b0),                               // (terminated)
		.reset_req_in7  (1'b0),                               // (terminated)
		.reset_in8      (1'b0),                               // (terminated)
		.reset_req_in8  (1'b0),                               // (terminated)
		.reset_in9      (1'b0),                               // (terminated)
		.reset_req_in9  (1'b0),                               // (terminated)
		.reset_in10     (1'b0),                               // (terminated)
		.reset_req_in10 (1'b0),                               // (terminated)
		.reset_in11     (1'b0),                               // (terminated)
		.reset_req_in11 (1'b0),                               // (terminated)
		.reset_in12     (1'b0),                               // (terminated)
		.reset_req_in12 (1'b0),                               // (terminated)
		.reset_in13     (1'b0),                               // (terminated)
		.reset_req_in13 (1'b0),                               // (terminated)
		.reset_in14     (1'b0),                               // (terminated)
		.reset_req_in14 (1'b0),                               // (terminated)
		.reset_in15     (1'b0),                               // (terminated)
		.reset_req_in15 (1'b0)                                // (terminated)
	);

endmodule
